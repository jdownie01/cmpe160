library ieee;
use ieee.std_logic_1164.all;


entity adder is
        port( a, b, cin         : in  STD_LOGIC;
              sum, cout         : out STD_LOGIC );
end adder;

architecture behaviorial of adder is
begin
	sum <=  (not a and not b and cin) or
                        (not a and b and not cin) or
                        (a and not b and not cin) or
                        (a and b and cin)after 8 ns;


    cout <= (not a and b and cin) or
                        (a and not b and cin) or
                        (a and b and not cin) or
                        (a and b and cin)after 8 ns;
end behaviorial;

